`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:43:18 02/10/2014 
// Design Name: 
// Module Name:    up_counter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module up_counter (sclr, clk, q);
  input sclr;
  input clk;
  output reg [19 : 0] q;
  
  always @(posedge clk)
  begin
	if(sclr)
		q <= 20'd0;
	else
		q <= q + 20'd1;
  end
  
endmodule
